library verilog;
use verilog.vl_types.all;
entity velocidade2_vlg_check_tst is
    port(
        c0              : in     vl_logic;
        c1              : in     vl_logic;
        c2              : in     vl_logic;
        c3              : in     vl_logic;
        c4              : in     vl_logic;
        c5              : in     vl_logic;
        c6              : in     vl_logic;
        c7              : in     vl_logic;
        clkout          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end velocidade2_vlg_check_tst;
