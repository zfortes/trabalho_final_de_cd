library verilog;
use verilog.vl_types.all;
entity velocidade2_vlg_vec_tst is
end velocidade2_vlg_vec_tst;
